-------------------------------------------------------------------------------
--
-- $Id: ttl_166-c.vhd,v 1.2 2005/10/10 22:12:38 arnim Exp $
--
-------------------------------------------------------------------------------

configuration ttl_166_rtl_c0 of ttl_166 is

  for rtl
  end for;

end ttl_166_rtl_c0;
