-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: prom_10_2-c.vhd,v 1.1 2005/11/15 23:51:54 arnim Exp $
--
-------------------------------------------------------------------------------

configuration prom_10_2_rtl_c0 of prom_10_2 is

  for rtl
  end for;

end prom_10_2_rtl_c0;
