-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: ladybug_addr_dec-c.vhd,v 1.2 2005/10/10 22:12:38 arnim Exp $
--
-------------------------------------------------------------------------------

configuration ladybug_addr_dec_rtl_c0 of ladybug_addr_dec is

  for rtl
  end for;

end ladybug_addr_dec_rtl_c0;
