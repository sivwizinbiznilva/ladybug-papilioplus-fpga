-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: rom_ram_dispatcher_16-c.vhd,v 1.1 2005/11/22 22:50:08 arnim Exp $
--
-------------------------------------------------------------------------------

configuration rom_ram_dispatcher_16_rtl_c0 of rom_ram_dispatcher_16 is

  for rtl
  end for;

end rom_ram_dispatcher_16_rtl_c0;
