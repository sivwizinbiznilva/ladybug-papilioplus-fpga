-------------------------------------------------------------------------------
--
-- $Id: pullup-c.vhd,v 1.1 2005/12/10 01:47:56 arnim Exp $
--
-------------------------------------------------------------------------------

configuration pullup_rtl_c0 of pullup is

  for rtl
  end for;

end pullup_rtl_c0;
