-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: ladybug_chute-c.vhd,v 1.2 2005/10/10 22:12:38 arnim Exp $
--
-------------------------------------------------------------------------------

configuration ladybug_chute_rtl_c0 of ladybug_chute is

  for rtl
  end for;

end ladybug_chute_rtl_c0;
