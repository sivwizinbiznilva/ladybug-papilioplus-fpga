-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: ladybug_por-altera-c.vhd,v 1.3 2005/11/07 21:56:12 arnim Exp $
--
-------------------------------------------------------------------------------

configuration ladybug_por_c0 of ladybug_por is

  for cyclone
  end for;

end ladybug_por_c0;
