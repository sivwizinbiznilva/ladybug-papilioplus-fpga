-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: ladybug_gpio-c.vhd,v 1.2 2005/10/10 22:12:38 arnim Exp $
--
-------------------------------------------------------------------------------

configuration ladybug_gpio_rtl_c0 of ladybug_gpio is

  for rtl
  end for;

end ladybug_gpio_rtl_c0;
