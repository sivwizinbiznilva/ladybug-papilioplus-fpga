-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: ladybug_clk-c.vhd,v 1.3 2005/10/28 21:17:32 arnim Exp $
--
-------------------------------------------------------------------------------

configuration ladybug_clk_rtl_c0 of ladybug_clk is

  for rtl
  end for;

end ladybug_clk_rtl_c0;
