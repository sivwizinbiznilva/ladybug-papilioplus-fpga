-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: prom_decrypt_l-c.vhd,v 1.1 2005/11/15 23:51:54 arnim Exp $
--
-------------------------------------------------------------------------------

configuration prom_decrypt_l_rtl_c0 of prom_decrypt_l is

  for rtl
  end for;

end prom_decrypt_l_rtl_c0;
