-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: generic_ram-c.vhd,v 1.1 2005/11/12 11:53:28 arnim Exp $
--
-------------------------------------------------------------------------------

configuration generic_ram_rtl_c0 of generic_ram is

  for rtl
  end for;

end generic_ram_rtl_c0;
