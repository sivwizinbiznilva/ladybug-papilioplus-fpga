-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: rom_dispatcher_8-c.vhd,v 1.1 2005/11/17 23:27:00 arnim Exp $
--
-------------------------------------------------------------------------------

configuration rom_dispatcher_8_rtl_c0 of rom_dispatcher_8 is

  for rtl
  end for;

end rom_dispatcher_8_rtl_c0;
