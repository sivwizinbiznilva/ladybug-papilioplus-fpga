-------------------------------------------------------------------------------
--
-- FPGA Lady Bug
--
-- $Id: prom_decrypt_u-c.vhd,v 1.1 2005/11/15 23:51:54 arnim Exp $
--
-------------------------------------------------------------------------------

configuration prom_decrypt_u_rtl_c0 of prom_decrypt_u is

  for rtl
  end for;

end prom_decrypt_u_rtl_c0;
